library ieee;
use ieee.std_logic_1164.ALL;
use ieee.numeric_std.ALL;


entity sm_ex3 is
	port(
	
	);
end sm_ex3;


architecture behavior of sm_ex3 is


end behavior;

